`timescale 1ns / 1ps

module Word_move(
    input [9:0] x_in,
    input [9:0] y_in,
    input [9:0] offset_x,
    input [9:0] offset_y,
    input [4:0] number,
    output logic display
    );
    
    logic [9:0] x, y;
    logic [0:62] word [31:0];
    
    assign x = x_in - offset_x;
    assign y = y_in - offset_y;
    
    assign word[0] = {
                            7'b0000000,
                            7'b0011100,
                            7'b0100010,
                            7'b0100110,
                            7'b0101010,
                            7'b0110010,
                            7'b0100010,
                            7'b0011100,
                            7'b0000000};
                            
    assign word[1] = {
                            7'b0000000,
                            7'b0001000,
                            7'b0011000,
                            7'b0001000,
                            7'b0001000,
                            7'b0001000,
                            7'b0001000,
                            7'b0011100,
                            7'b0000000};
                            
    assign word[2] = {
                            7'b0000000,
                            7'b0011100,
                            7'b0100010,
                            7'b0000010,
                            7'b0000100,
                            7'b0001000,
                            7'b0010000,
                            7'b0111110,
                            7'b0000000};
                            
    assign word[3] = {
                            7'b0000000,
                            7'b0111110,
                            7'b0000100,
                            7'b0001000,
                            7'b0000100,
                            7'b0000010,
                            7'b0100010,
                            7'b0011100,
                            7'b0000000};
                            
    assign word[4] = {
                            7'b0000000,
                            7'b0000100,
                            7'b0001100,
                            7'b0010100,
                            7'b0100100,
                            7'b0111110,
                            7'b0000100,
                            7'b0000100,
                            7'b0000000};
                               
    assign word[5] = {
                            7'b0000000,
                            7'b0111110,
                            7'b0100000,
                            7'b0111100,
                            7'b0000010,
                            7'b0000010,
                            7'b0100010,
                            7'b0011100,
                            7'b0000000};
                            
    assign word[6] = {
                            7'b0000000,
                            7'b0001100,
                            7'b0010000,
                            7'b0100000,
                            7'b0111100,
                            7'b0100010,
                            7'b0100010,
                            7'b0011100,
                            7'b0000000};
                            
    assign word[7] = {
                            7'b0000000,
                            7'b0111110,
                            7'b0000010,
                            7'b0000100,
                            7'b0001000,
                            7'b0010000,
                            7'b0010000,
                            7'b0010000,
                            7'b0000000};
                            
    assign word[8] = {
                            7'b0000000,
                            7'b0011100,
                            7'b0100010,
                            7'b0100010,
                            7'b0011100,
                            7'b0100010,
                            7'b0100010,
                            7'b0011100,
                            7'b0000000};
                            
    assign word[9] = {
                            7'b0000000,
                            7'b0011100,
                            7'b0100010,
                            7'b0100010,
                            7'b0011110,
                            7'b0000010,
                            7'b0000100,
                            7'b0011000,
                            7'b0000000};
                            
    assign word[10] = {
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0011000,
                            7'b0011000,
                            7'b0000000};
                                                                              
    assign word[11] = {
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0110100,
                            7'b0101010,
                            7'b0101010,
                            7'b0100010,
                            7'b0100010,
                            7'b0000000};
                                                                              
    assign word[12] = {
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0100010,
                            7'b0100010,
                            7'b0100010,
                            7'b0100110,
                            7'b0111010,
                            7'b0100000};
                                                                              
    assign word[13] = {
                            7'b0000000,
                            7'b0100010,
                            7'b0100010,
                            7'b0100010,
                            7'b0100010,
                            7'b0100010,
                            7'b0010100,
                            7'b0001000,
                            7'b0000000};
                                                                              
    assign word[14] = {
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0111110,
                            7'b0000000,
                            7'b0101010,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000};

                                                                              
    assign word[15] = {
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0010000,
                            7'b0101010,
                            7'b0000100,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000};                                                      
                                                                              
    assign word[16] = {
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000};   
                                                                              
    assign word[17] = {
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0111110,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000,
                            7'b0000000};
 
     assign word[18] = {
                            7'b0000000,
                            7'b0001110,
                            7'b0001000,
                            7'b0001000,
                            7'b0011100,
                            7'b0111110,
                            7'b0001000,
                            7'b0111000,
                            7'b0000000};
                                                                                                                                                                                                                                                            
    assign display = (x <= 6 & y <= 8)? word[number][y*7+x] : 0;
    
endmodule
